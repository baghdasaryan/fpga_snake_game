----------------------------------------------------------------------------------
-- Engineer: Georgi Baghdasaryan, UID: 603 875 284
-- 
-- Create Date:    05/24/2013 
-- Project Name:   Lab 6: Final Project (Snake Game)
-- Target Devices: Spartan 3 Board
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity display is
  port(clk50_in  : in STD_LOGIC;
       reset_in  : in STD_LOGIC;
		 win_in    : in STD_LOGIC;
       appleX_in : in integer range 0 to 630;
       appleY_in : in integer range 0 to 470;
       move_in   : in STD_LOGIC_VECTOR(1 downto 0);
       rgb_out   : out STD_LOGIC_VECTOR(2 downto 0);
       hs_out    : out STD_LOGIC;
       vs_out    : out STD_LOGIC;
		 game_out  : out STD_LOGIC;
		 score_out : out STD_LOGIC);
end display ;

architecture Behavioral of display is

signal clk25     : STD_LOGIC;
signal hcounter  : integer range 0 to 800;
signal vcounter  : integer range 0 to 521;

signal speed     : integer range 0 to 31 := 1;
signal gameOver  : STD_LOGIC := '0';
signal refresh   : STD_LOGIC := '0';

-- Location
type POS is array (29 downto 0, 1 downto 0) of integer;
type TEMP is array (1 downto 0) of integer;
signal my_pos : POS;
signal apple  : TEMP := (appleY_in,appleX_in);

-- Object colors
constant border_color: STD_LOGIC_VECTOR(2 downto 0) := "001";
constant snake_color	: STD_LOGIC_VECTOR(2 downto 0) := "010";
constant apple_color	: STD_LOGIC_VECTOR(2 downto 0) := "100";
constant back_color	: STD_LOGIC_VECTOR(2 downto 0) := "000";

-- Text
type GO is array (19 downto 0) of STD_LOGIC_VECTOR(221 downto 0);
constant gameOverText : GO := (
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110",
"000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
"000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
"001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
"011111110000000111111000000011111111111110000000000011111110000111111100000000000011111111111100000000000000000001111111100011111111000001111111000000000001111111000000000111111111111000000000111110001111111110000000011111",
"111111100000000000000000000011111111111111000000001111111111001111111111000000001111111111111111000000000000000001111111000001111111000000111111100000000011111110000000011111111111111110000000111111111111111111000000011111",
"111111100000000000000000000011111111111111100000011111111111111111111111100000011111111111111111110000000000000001111111000001111111000000011111110000000111111100000000111111111111111111100000111111111111111111100000011111",
"111111100001111111111000000000000000011111100000011111111111111111111111100000111111110000011111110000000000000001111111000001111111000000001111111000001111111000000001111111100000111111100000111111111111111111110000011111",
"111111100001111111111000000000111111111111100000011111111111111111111111100000111111111111111111110000000000000001111111000001111111000000000111111100011111110000000001111111111111111111100000011111110000011111110000011111",
"111111100001111111111000000011111111111111100000011111100011111100011111100000111111111111111111100000000000000001111111000001111111000000000011111110111111100000000001111111111111111111000000011111110000011111110000011111",
"111111100000000111111000000111111111111111100000011111100011111100011111100000111111111111111111000000000000000001111111000001111111000000000001111111111111000000000001111111111111111110000000011111110000000000000000011111",
"011111110000000111111000001111110000111111100000011111100011111100011111100000111111111000000000000000000000000001111111100011111111000000000000111111111110000000000001111111110000000000000000011111110000000000000000001110",
"001111111111111111111000001111110000111111100000011111100011111100011111100000111111111100000000000000000000000001111111111111111111000000000000011111111100000000000001111111111000000000000000011111110000000000000000000000",
"000111111111111111111000001111111111111111100000011111100011111100011111100000011111111111111111000000000000000000111111111111111110000000000000001111111000000000000000111111111111111110000000011111110000000000000000001110",
"000001111111111111111000000111111111111111110000011111100011111100011111100000001111111111111111000000000000000000001111111111111000000000000000000111110000000000000000011111111111111110000000011111110000000000000000011111",
"000000001111110001111000000011111111110011110000011111100011111100011111100000000011111111111111000000000000000000000011111111100000000000000000000011100000000000000000000111111111111110000000011111110000000000000000001110",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");

type YO is array (19 downto 0) of STD_LOGIC_VECTOR(178 downto 0);
constant youWonText : YO := (
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"11111110000000111111100000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000111111110000000000000000000000000000000000000000000000000001110",
"11111110000000111111100000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000111111110000000000000000000000000000000000000000000000000011111",
"11111110000000111111100000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000111111110000000000000000000000000000000000000000000000000011111",
"11111111000001111111100000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000111111110000000000000000000000000000000000000000000000000011111",
"11111111100011111111100000000111111111110000000011111100001111110000000000000000001111111000000000001111100000000000111111100000000011111111111000000001111001111111100000000011111",
"00011111110111111100000000011111111111111100000011111100001111110000000000000000000111111100000000011111110000000001111111000000001111111111111110000001111111111111111000000011111",
"00001111111111111000000000111111111111111110000011111100001111110000000000000000000011111110000000111111111000000011111110000000011111111111111111000001111111111111111100000011111",
"00000111111111110000000000111111111111111110000011111100001111110000000000000000000001111111000001111111111100000111111100000000011111111111111111000001111111111111111110000011111",
"00000011111111100000000000111111000001111110000011111100001111110000000000000000000000111111100011111111111110001111111000000000011111100000111111000000011111111111111110000011111",
"00000001111111000000000000111111000001111110000011111100001111110000000000000000000000011111110111111101111111011111110000000000011111100000111111000000011111100001111110000011111",
"00000001111111000000000000111111000001111110000011111100001111110000000000000000000000001111111111111000111111111111100000000000011111100000111111000000011111100001111110000011111",
"00000001111111000000000000111111000001111110000011111111111111110000000000000000000000000111111111110000011111111111000000000000011111100000111111000000011111100001111110000001110",
"00000001111111000000000000111111111111111110000011111111111111111100000000000000000000000011111111100000001111111110000000000000011111111111111111000000011111100001111110000000000",
"00001111111111111000000000111111111111111110000001111111111111111100000000000000000000000001111111000000000111111100000000000000011111111111111111000000011111100001111110000001110",
"00001111111111111000000000011111111111111100000000111111111111111100000000000000000000000000111110000000000011111000000000000000001111111111111110000000011111100001111110000011111",
"00001111111111111000000000000111111111110000000000001111111100111100000000000000000000000000011100000000000001110000000000000000000011111111111000000000011111100001111110000001110",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");


begin
	
	-- Generate a 25Mhz clock
	process(clk50_in)
	begin
	  if clk50_in'event and clk50_in='1' then
		 clk25 <= not clk25;
	  end if;
	end process;

	-- Horizontal and vertical clocks
	process(clk25)
	begin
		if clk25'event and clk25 = '1' then
			if hcounter = 800 then
				hcounter <= 0;
				if vcounter = 521 then
					vcounter <= 0;
					refresh <= refresh xor '1';
				else
					vcounter <= vcounter + 1;
				end if;
			else
				hcounter <= hcounter + 1;
			end if;
		end if;
	end process;
	
	process (clk25, hcounter, vcounter, gameOver, win_in)
		variable x: integer range 0 to 639;
		variable y: integer range 0 to 479;
	begin
		-- hcounter counts from 0 to 799
		-- vcounter counts from 0 to 520
		-- x coordinate: 0 - 639 (x = hcounter - 144, i.e., hcounter -Tpw-Tbp)
		-- y coordinate: 0 - 479 (y = vcounter - 31, i.e., vcounter-Tpw-Tbp)
		x := hcounter - 144;
		y := vcounter - 31;
		if clk25'event and clk25 = '1' then
			
			if x < 640 and y < 480 and gameOver = '0' and win_in = '0' then
				-- Display borders, snake, apples, and background				
				if y <= 10 or y >= 470 or x >= 630 or x <= 10 then
					rgb_out <= border_color;
				elsif (x >= apple(0) - 5 and x <= apple(0) + 5 and y >= apple(1) - 5 and y <= apple(1) + 5) and reset_in = '0' then
					rgb_out <= apple_color;
				else
					rgb_out <= back_color;
				end if;
				for i in 0 to 5 loop
					if (x >= (integer(my_pos(i,0) - 5)) and x <= (integer(my_pos(i,0) + 5)) and y >= (integer(my_pos(i,1) - 5)) and y <= (integer(my_pos(i,1) + 5))) then  -- add offsets
						rgb_out <= snake_color;
					end if;
				end loop;
			elsif gameOver = '1' then
				if x >= 208 and x <= 430 and y >= 129 and y <= 350 then
					if gameOverText(19-(y-129))(221-(x-208)) = '1' then
						rgb_out <= apple_color;
					else
						rgb_out <= back_color;
					end if;
				end if;
			elsif win_in = '1' then
				if x >= 230 and x <= 410 and y >= 129 and y <= 350 then
					if youWonText(19-(y-129))(178-(x-230)) = '1' then
						rgb_out <= snake_color;
					else
						rgb_out <= back_color;
					end if;
				end if;
			else
				-- If not traced, set it to "black" color
				rgb_out <= back_color;
			end if;
			
			-- Set horizontal and vertical synchronizations.
			if hcounter < 96 then
				hs_out <= '0';
			else
				hs_out <= '1';
			end if;
			if vcounter < 2 then
				vs_out <= '0';
			else
				vs_out <= '1';
			end if;
			
	  end if;
	end process;

	-- Update snake's location
	process(refresh, reset_in, move_in, gameOver)
	begin
		if refresh'event and refresh = '1' then
			
			for i in 1 to 5 loop
--				if ((integer(my_pos(0,0) + 5) >= integer(my_pos(i,0) - 5)) and (integer(my_pos(0,0) + 5) <= integer(my_pos(i,0) + 5))) or ((integer(my_pos(0,0) - 5) >= integer(my_pos(i,0) - 5)) and (integer(my_pos(0,0) - 5) <= integer(my_pos(i,0) + 5))) or ((integer(my_pos(0,1) - 5) >= integer(my_pos(i,1) - 5)) and (integer(my_pos(0,1) - 5) <= integer(my_pos(i,0) + 5)))or ((integer(my_pos(0,1) + 5) >= integer(my_pos(i,1) - 5)) and (integer(my_pos(0,1) + 5) <= integer(my_pos(i,0) + 5))) then
--					gameOver <= '1';
--				end if;
				my_pos(i,0) <= my_pos(i-1,0);
				my_pos(i,1) <= my_pos(i-1,1);
			end loop;
			
			if reset_in = '1' then
				for i in 0 to 5 loop
					my_pos(i,0) <= 320;
					my_pos(i,1) <= 240;
				end loop;
				apple <= (appleY_in,appleX_in);
				speed <= 1;
				gameOver <= '0';
			elsif (my_pos(0,0) + 5) >= 630 or (my_pos(0,0) - 5) <= 10 or (my_pos(0,1) + 5) >= 470 or (my_pos(0,1) - 5) <= 10 then
				gameOver <= '1';
			elsif move_in = "00" then
				my_pos(0,0) <= my_pos(0,0) + speed;
			elsif move_in = "01" then
				my_pos(0,0) <= my_pos(0,0) - speed;
			elsif move_in = "10" then
				my_pos(0,1) <= my_pos(0,1) - speed;
			else
				my_pos(0,1) <= my_pos(0,1) + speed;
			end if;
			
			if (((my_pos(0,0)-5 >= apple(0)-5) and (my_pos(0,0)-5 <= apple(0)+5)) or ((my_pos(0,0)+5 >= apple(0)-5) and (my_pos(0,0)+5 <= apple(0)+5))) and 
				(((my_pos(0,1)-5 >= apple(1)-5) and (my_pos(0,1)-5 <= apple(1)+5)) or ((my_pos(0,1)+5 >= apple(1)-5) and (my_pos(0,1)+5 <= apple(1)+5))) then
				score_out <= '1';
				apple <= (appleY_in,appleX_in);
				speed <= speed + 1;
			else
				score_out <= '0';
			end if;
			
		end if;
	end process;
	
	-- Set game output
	process(gameOver)
	begin
		if gameOver = '1' then
			game_out <= '1';
		else
			game_out <= '0';
		end if;
	end process;
	
end Behavioral;

